.title KiCad schematic
P1 NC_01 NC_02 NC_03 /SLTSL NC_04 NC_05 /WAIT /INT /M1 /BUSDIR /IORQ /MREQ /WR /RD NC_06 NC_07 /A9 /A15 /A11 /A10 /A7 /A6 /A12 /A8 /A14 /A13 /A1 /A0 /A3 /A2 /A5 /A4 /D1 /D0 /D3 /D2 /D5 /D4 /D7 /D6 GND /CLK GND Net-_P1-Pad44_ +5V Net-_P1-Pad44_ +5V NC_08 /SOUNDIN NC_09 CONN_02X25
U5 +5V /DAT_DIR /D1 /D0 /D3 /D2 /D5 /D4 /D7 /D6 GND GND GND /RD6 /RD7 /RD4 /RD5 /RD2 /RD3 /RD0 /RD1 /DAT_EN +3V3 +3V3 LVC4245
U4 GND /CLK /RC19 /M1 /RC26 /WR /RC17 /RD NC_10 GND NC_11 /RC20 /SLTSL /RC27 /MREQ /RC21 /IORQ NC_12 GND +3V3 74HC244
J1 +3V3 +5V /RD2 +5V /RD3 GND /RD4 NC_13 GND NC_14 /RC17 /RC18 /RC27 GND /ADDR /RC23 +3V3 /RC24 NC_15 GND NC_16 /DAT_DIR NC_17 NC_18 GND /RD7 /RD0 /RD1 /RD5 GND /RD6 NC_19 NC_20 GND /RC19 /DAT_EN /RC26 /RC20 GND /RC21 RPi_GPIO
D1 /DAT_EN /SLTSL /DAT_DIR Net-_D1-Pad4_ Net-_D1-Pad5_ Net-_D1-Pad6_ LED_RGB
R1 Net-_D1-Pad6_ +3V3 R
R2 Net-_D1-Pad5_ +3V3 R
R3 Net-_D1-Pad4_ +3V3 R
U3 /CWAIT /WAIT /RC23 /INT /DAT_DIR /BUSDIR 74LS07
J2 /RD2 /RD3 +3V3 GND Conn_01x04
C2 GND Net-_C1-Pad1_ C
C1 Net-_C1-Pad1_ /SOUNDIN CP
R4 Net-_C1-Pad1_ /RC18 R
R5 GND Net-_C1-Pad1_ R
U1 /ADDR /A8 NC_21 /A9 NC_22 /A10 NC_23 /A11 NC_24 GND /A15 NC_25 /A14 NC_26 /A13 NC_27 /A12 NC_28 /ADDR +3V3 74HC244
U2 /ADDR /A6 /RD2 /A7 /RD3 /A4 /RD0 /A5 /RD1 GND /A1 /RD5 /A0 /RD4 /A3 /RD7 /A2 /RD6 /ADDR +3V3 74HC244
U6 /IORQ /MREQ Net-_U6-Pad3_ Net-_U6-Pad3_ /RC24 /CWAIT 74HC00
.end
