// plltest.v

// Generated using ACDS version 13.1 162 at 2016.03.02.01:21:33

`timescale 1 ps / 1 ps
module plltest (
		input  wire  clk_clk,       //       clk.clk
		input  wire  reset_reset_n, //     reset.reset_n
		output wire  clk_0_clk_clk  // clk_0_clk.clk
	);

	assign clk_0_clk_clk = clk_clk;

endmodule
